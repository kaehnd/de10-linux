// DE10_Linux.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module DE10_Linux (
		input  wire        clk_clk,                   //   clk.clk
		input  wire        reset_reset_n,             // reset.reset_n
		output wire [12:0] sdram_sdram_addr,          // sdram.sdram_addr
		output wire [1:0]  sdram_sdram_ba,            //      .sdram_ba
		output wire        sdram_new_signal,          //      .new_signal
		output wire        sdram_sdram_chipselect_n,  //      .sdram_chipselect_n
		inout  wire [15:0] sdram_sdram_dq,            //      .sdram_dq
		output wire [1:0]  sdram_sdram_dqm,           //      .sdram_dqm
		output wire        sdram_sdram_ras_n,         //      .sdram_ras_n
		output wire        sdram_sdram_writeenable_n, //      .sdram_writeenable_n
		output wire        sdram_sdram_cke            //      .sdram_cke
	);

	wire         altpll_0_c0_clk;                                                // altpll_0:c0 -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, mm_interconnect_2:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, onchip_memory2_0:clk2, rst_controller_002:clk, rst_controller_003:clk]
	wire         altpll_0_c1_clk;                                                // altpll_0:c1 -> [de10_lite_sdram_0:clk, mm_interconnect_0:altpll_0_c1_clk, rst_controller_001:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                              // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                           // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                           // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                               // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                            // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                  // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                         // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                 // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                             // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                       // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                        // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                           // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                  // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_de10_lite_sdram_0_avalon_slave_chipselect;    // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_chipselect -> de10_lite_sdram_0:az_cs
	wire  [15:0] mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdata;      // de10_lite_sdram_0:za_data -> mm_interconnect_0:de10_lite_sdram_0_avalon_slave_readdata
	wire         mm_interconnect_0_de10_lite_sdram_0_avalon_slave_waitrequest;   // de10_lite_sdram_0:za_waitrequest -> mm_interconnect_0:de10_lite_sdram_0_avalon_slave_waitrequest
	wire  [24:0] mm_interconnect_0_de10_lite_sdram_0_avalon_slave_address;       // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_address -> de10_lite_sdram_0:az_addr
	wire         mm_interconnect_0_de10_lite_sdram_0_avalon_slave_read;          // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_read -> de10_lite_sdram_0:az_rd_n
	wire   [1:0] mm_interconnect_0_de10_lite_sdram_0_avalon_slave_byteenable;    // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_byteenable -> de10_lite_sdram_0:az_be_n
	wire         mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdatavalid; // de10_lite_sdram_0:za_valid -> mm_interconnect_0:de10_lite_sdram_0_avalon_slave_readdatavalid
	wire         mm_interconnect_0_de10_lite_sdram_0_avalon_slave_write;         // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_write -> de10_lite_sdram_0:az_wr_n
	wire  [15:0] mm_interconnect_0_de10_lite_sdram_0_avalon_slave_writedata;     // mm_interconnect_0:de10_lite_sdram_0_avalon_slave_writedata -> de10_lite_sdram_0:az_data
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;        // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;     // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                  // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                   // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                      // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                     // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                 // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] nios2_gen2_0_tightly_coupled_data_master_0_readdata;            // mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_readdata -> nios2_gen2_0:dtcm0_readdata
	wire  [15:0] nios2_gen2_0_tightly_coupled_data_master_0_address;             // nios2_gen2_0:dtcm0_address -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_address
	wire         nios2_gen2_0_tightly_coupled_data_master_0_read;                // nios2_gen2_0:dtcm0_read -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_read
	wire   [3:0] nios2_gen2_0_tightly_coupled_data_master_0_byteenable;          // nios2_gen2_0:dtcm0_byteenable -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_byteenable
	wire         nios2_gen2_0_tightly_coupled_data_master_0_write;               // nios2_gen2_0:dtcm0_write -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_write
	wire  [31:0] nios2_gen2_0_tightly_coupled_data_master_0_writedata;           // nios2_gen2_0:dtcm0_writedata -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_writedata
	wire         nios2_gen2_0_tightly_coupled_data_master_0_clken;               // nios2_gen2_0:dtcm0_clken -> mm_interconnect_1:nios2_gen2_0_tightly_coupled_data_master_0_clken
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;               // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;                 // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_1_onchip_memory2_0_s1_address;                  // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;               // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;                    // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;                // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;                    // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] nios2_gen2_0_tightly_coupled_instruction_master_0_readdata;     // mm_interconnect_2:nios2_gen2_0_tightly_coupled_instruction_master_0_readdata -> nios2_gen2_0:itcm0_readdata
	wire  [15:0] nios2_gen2_0_tightly_coupled_instruction_master_0_address;      // nios2_gen2_0:itcm0_address -> mm_interconnect_2:nios2_gen2_0_tightly_coupled_instruction_master_0_address
	wire         nios2_gen2_0_tightly_coupled_instruction_master_0_read;         // nios2_gen2_0:itcm0_read -> mm_interconnect_2:nios2_gen2_0_tightly_coupled_instruction_master_0_read
	wire         nios2_gen2_0_tightly_coupled_instruction_master_0_clken;        // nios2_gen2_0:itcm0_clken -> mm_interconnect_2:nios2_gen2_0_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_2_onchip_memory2_0_s2_chipselect;               // mm_interconnect_2:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_2_onchip_memory2_0_s2_readdata;                 // onchip_memory2_0:readdata2 -> mm_interconnect_2:onchip_memory2_0_s2_readdata
	wire  [13:0] mm_interconnect_2_onchip_memory2_0_s2_address;                  // mm_interconnect_2:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_2_onchip_memory2_0_s2_byteenable;               // mm_interconnect_2:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_2_onchip_memory2_0_s2_write;                    // mm_interconnect_2:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_2_onchip_memory2_0_s2_writedata;                // mm_interconnect_2:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_2_onchip_memory2_0_s2_clken;                    // mm_interconnect_2:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire         irq_mapper_receiver0_irq;                                       // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                           // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [de10_lite_sdram_0:reset_n, mm_interconnect_0:de10_lite_sdram_0_reset_n_reset_bridge_in_reset_reset]
	wire         nios2_gen2_0_debug_reset_request_reset;                         // nios2_gen2_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                             // rst_controller_002:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                         // rst_controller_002:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                             // rst_controller_003:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset2, rst_translator_001:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                         // rst_controller_003:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator_001:reset_req_in]

	DE10_Linux_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (altpll_0_c1_clk),                                //                    c1.clk
		.areset             (),                                               //        areset_conduit.export
		.locked             (),                                               //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	DE10_LITE_Qsys_sdram de10_lite_sdram_0 (
		.clk            (altpll_0_c1_clk),                                                //          clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                            //      reset_n.reset_n
		.az_addr        (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_address),       // avalon_slave.address
		.az_be_n        (~mm_interconnect_0_de10_lite_sdram_0_avalon_slave_byteenable),   //             .byteenable_n
		.az_cs          (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_chipselect),    //             .chipselect
		.az_rd_n        (~mm_interconnect_0_de10_lite_sdram_0_avalon_slave_read),         //             .read_n
		.az_wr_n        (~mm_interconnect_0_de10_lite_sdram_0_avalon_slave_write),        //             .write_n
		.az_data        (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_writedata),     //             .writedata
		.za_data        (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdata),      //             .readdata
		.za_waitrequest (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_waitrequest),   //             .waitrequest
		.za_valid       (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdatavalid), //             .readdatavalid
		.zs_addr        (sdram_sdram_addr),                                               //        sdram.sdram_addr
		.zs_ba          (sdram_sdram_ba),                                                 //             .sdram_ba
		.zs_cas_n       (sdram_new_signal),                                               //             .new_signal
		.zs_cs_n        (sdram_sdram_chipselect_n),                                       //             .sdram_chipselect_n
		.zs_dq          (sdram_sdram_dq),                                                 //             .sdram_dq
		.zs_dqm         (sdram_sdram_dqm),                                                //             .sdram_dqm
		.zs_ras_n       (sdram_sdram_ras_n),                                              //             .sdram_ras_n
		.zs_we_n        (sdram_sdram_writeenable_n),                                      //             .sdram_writeenable_n
		.zs_cke         (sdram_sdram_cke)                                                 //             .sdram_cke
	);

	DE10_Linux_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	DE10_Linux_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                                  clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                        //                                reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),                     //                                     .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //                          data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                                     .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                                     .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                                     .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                                     .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                                     .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                                     .readdatavalid
		.dtcm0_readdata                      (nios2_gen2_0_tightly_coupled_data_master_0_readdata),        //        tightly_coupled_data_master_0.readdata
		.dtcm0_address                       (nios2_gen2_0_tightly_coupled_data_master_0_address),         //                                     .address
		.dtcm0_read                          (nios2_gen2_0_tightly_coupled_data_master_0_read),            //                                     .read
		.dtcm0_clken                         (nios2_gen2_0_tightly_coupled_data_master_0_clken),           //                                     .clken
		.dtcm0_write                         (nios2_gen2_0_tightly_coupled_data_master_0_write),           //                                     .write
		.dtcm0_writedata                     (nios2_gen2_0_tightly_coupled_data_master_0_writedata),       //                                     .writedata
		.dtcm0_byteenable                    (nios2_gen2_0_tightly_coupled_data_master_0_byteenable),      //                                     .byteenable
		.itcm0_readdata                      (nios2_gen2_0_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (nios2_gen2_0_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (nios2_gen2_0_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (nios2_gen2_0_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                     .writedata
		.dummy_ci_port                       ()                                                            //            custom_instruction_master.readra
	);

	DE10_Linux_onchip_memory2_0 onchip_memory2_0 (
		.clk         (altpll_0_c0_clk),                                  //   clk1.clk
		.address     (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_002_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_002_reset_out_reset_req),           //       .reset_req
		.address2    (mm_interconnect_2_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk2        (altpll_0_c0_clk),                                  //   clk2.clk
		.reset2      (rst_controller_003_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_003_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	DE10_Linux_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                                //                                          altpll_0_c0.clk
		.altpll_0_c1_clk                                            (altpll_0_c1_clk),                                                //                                          altpll_0_c1.clk
		.clk_0_clk_clk                                              (clk_clk),                                                        //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.de10_lite_sdram_0_reset_n_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                             //      de10_lite_sdram_0_reset_n_reset_bridge_in_reset.reset
		.jtag_uart_0_reset_reset_bridge_in_reset_reset              (rst_controller_002_reset_out_reset),                             //              jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                             //             nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                               //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                           //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                            //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                  //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                              //                                                     .readdata
		.nios2_gen2_0_data_master_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                         //                                                     .readdatavalid
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                 //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                             //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                           //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                        //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                    //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                           //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                       //                                                     .readdata
		.nios2_gen2_0_instruction_master_readdatavalid              (nios2_gen2_0_instruction_master_readdatavalid),                  //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                   //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                     //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                      //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                  //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                 //                                                     .writedata
		.de10_lite_sdram_0_avalon_slave_address                     (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_address),       //                       de10_lite_sdram_0_avalon_slave.address
		.de10_lite_sdram_0_avalon_slave_write                       (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_write),         //                                                     .write
		.de10_lite_sdram_0_avalon_slave_read                        (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_read),          //                                                     .read
		.de10_lite_sdram_0_avalon_slave_readdata                    (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdata),      //                                                     .readdata
		.de10_lite_sdram_0_avalon_slave_writedata                   (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_writedata),     //                                                     .writedata
		.de10_lite_sdram_0_avalon_slave_byteenable                  (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_byteenable),    //                                                     .byteenable
		.de10_lite_sdram_0_avalon_slave_readdatavalid               (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_readdatavalid), //                                                     .readdatavalid
		.de10_lite_sdram_0_avalon_slave_waitrequest                 (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_waitrequest),   //                                                     .waitrequest
		.de10_lite_sdram_0_avalon_slave_chipselect                  (mm_interconnect_0_de10_lite_sdram_0_avalon_slave_chipselect),    //                                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),         //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),           //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),            //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),        //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),       //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),      //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),     //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess)      //                                                     .debugaccess
	);

	DE10_Linux_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                                       (altpll_0_c0_clk),                                       //                                   altpll_0_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset        (rst_controller_003_reset_out_reset),                    //      nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset   (rst_controller_002_reset_out_reset),                    // onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.nios2_gen2_0_tightly_coupled_data_master_0_address    (nios2_gen2_0_tightly_coupled_data_master_0_address),    //    nios2_gen2_0_tightly_coupled_data_master_0.address
		.nios2_gen2_0_tightly_coupled_data_master_0_byteenable (nios2_gen2_0_tightly_coupled_data_master_0_byteenable), //                                              .byteenable
		.nios2_gen2_0_tightly_coupled_data_master_0_read       (nios2_gen2_0_tightly_coupled_data_master_0_read),       //                                              .read
		.nios2_gen2_0_tightly_coupled_data_master_0_readdata   (nios2_gen2_0_tightly_coupled_data_master_0_readdata),   //                                              .readdata
		.nios2_gen2_0_tightly_coupled_data_master_0_write      (nios2_gen2_0_tightly_coupled_data_master_0_write),      //                                              .write
		.nios2_gen2_0_tightly_coupled_data_master_0_writedata  (nios2_gen2_0_tightly_coupled_data_master_0_writedata),  //                                              .writedata
		.nios2_gen2_0_tightly_coupled_data_master_0_clken      (nios2_gen2_0_tightly_coupled_data_master_0_clken),      //                                              .clken
		.onchip_memory2_0_s1_address                           (mm_interconnect_1_onchip_memory2_0_s1_address),         //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                             (mm_interconnect_1_onchip_memory2_0_s1_write),           //                                              .write
		.onchip_memory2_0_s1_readdata                          (mm_interconnect_1_onchip_memory2_0_s1_readdata),        //                                              .readdata
		.onchip_memory2_0_s1_writedata                         (mm_interconnect_1_onchip_memory2_0_s1_writedata),       //                                              .writedata
		.onchip_memory2_0_s1_byteenable                        (mm_interconnect_1_onchip_memory2_0_s1_byteenable),      //                                              .byteenable
		.onchip_memory2_0_s1_chipselect                        (mm_interconnect_1_onchip_memory2_0_s1_chipselect),      //                                              .chipselect
		.onchip_memory2_0_s1_clken                             (mm_interconnect_1_onchip_memory2_0_s1_clken)            //                                              .clken
	);

	DE10_Linux_mm_interconnect_2 mm_interconnect_2 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                            //                                       altpll_0_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                         //          nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_tightly_coupled_instruction_master_0_address  (nios2_gen2_0_tightly_coupled_instruction_master_0_address),  // nios2_gen2_0_tightly_coupled_instruction_master_0.address
		.nios2_gen2_0_tightly_coupled_instruction_master_0_read     (nios2_gen2_0_tightly_coupled_instruction_master_0_read),     //                                                  .read
		.nios2_gen2_0_tightly_coupled_instruction_master_0_readdata (nios2_gen2_0_tightly_coupled_instruction_master_0_readdata), //                                                  .readdata
		.nios2_gen2_0_tightly_coupled_instruction_master_0_clken    (nios2_gen2_0_tightly_coupled_instruction_master_0_clken),    //                                                  .clken
		.onchip_memory2_0_s2_address                                (mm_interconnect_2_onchip_memory2_0_s2_address),              //                               onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                                  (mm_interconnect_2_onchip_memory2_0_s2_write),                //                                                  .write
		.onchip_memory2_0_s2_readdata                               (mm_interconnect_2_onchip_memory2_0_s2_readdata),             //                                                  .readdata
		.onchip_memory2_0_s2_writedata                              (mm_interconnect_2_onchip_memory2_0_s2_writedata),            //                                                  .writedata
		.onchip_memory2_0_s2_byteenable                             (mm_interconnect_2_onchip_memory2_0_s2_byteenable),           //                                                  .byteenable
		.onchip_memory2_0_s2_chipselect                             (mm_interconnect_2_onchip_memory2_0_s2_chipselect),           //                                                  .chipselect
		.onchip_memory2_0_s2_clken                                  (mm_interconnect_2_onchip_memory2_0_s2_clken)                 //                                                  .clken
	);

	DE10_Linux_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c1_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
